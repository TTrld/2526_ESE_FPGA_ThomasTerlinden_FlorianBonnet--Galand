library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library pll;
use pll.all;

entity telecran is
    port (
        -- FPGA
        i_clk_50 : in std_logic;

        -- HDMI
        io_hdmi_i2c_scl : inout std_logic;
        io_hdmi_i2c_sda : inout std_logic;
        o_hdmi_tx_clk   : out std_logic;
        o_hdmi_tx_d     : out std_logic_vector(23 downto 0);
        o_hdmi_tx_de    : out std_logic;
        o_hdmi_tx_hs    : out std_logic;
        i_hdmi_tx_int   : in std_logic;
        o_hdmi_tx_vs    : out std_logic;

        -- KEYs
        i_rst_n : in std_logic;

        -- LEDs
        o_leds : out std_logic_vector(9 downto 0);
        o_de10_leds : out std_logic_vector(7 downto 0);

        -- Coder
        i_left_ch_a : in std_logic;--Axe X
        i_left_ch_b : in std_logic;
        i_left_pb   : in std_logic;
        i_right_ch_a : in std_logic;--Axe Y
        i_right_ch_b : in std_logic;
        i_right_pb   : in std_logic
    );
end entity telecran;

architecture rtl of telecran is

    component I2C_HDMI_Config 
        port (
            iCLK : in std_logic;
            iRST_N : in std_logic;
            I2C_SCLK : out std_logic;
            I2C_SDAT : inout std_logic;
            HDMI_TX_INT  : in std_logic
        );
    end component;
    
    component pll 
        port (
            refclk : in std_logic;
            rst : in std_logic;
            outclk_0 : out std_logic;
            locked : out std_logic
        );
    end component;

    constant h_res : natural := 720;
    constant v_res : natural := 480;

    signal s_clk_27 : std_logic;
    signal s_rst_n : std_logic; -- holds reset as long as pll is not locked
	 
	 -- Signaux pour récupérer la position de balayage du contrôleur HDMI
    signal s_scan_x : unsigned(11 downto 0);
    signal s_scan_y : unsigned(11 downto 0);
    signal s_de     : std_logic; -- Data Enable interne

	 -- Signaux Position Curseur (sorties des instances encodeurs)
    signal s_pos_x  : integer range 0 to h_res-1;
    signal s_pos_y  : integer range 0 to v_res-1;

	 -- On change la taille des vecteurs de données mémoire à 1 bit
    signal s_pixel_data : std_logic_vector(0 downto 0); 
    signal s_data_a     : std_logic_vector(0 downto 0);
    
    signal s_we_a       : std_logic;
    signal s_addr_a     : natural range 0 to h_res*v_res-1;

begin
    o_leds <= (others => '0');
    o_de10_leds <= (others => '0');
    
    -- Frequency for HDMI is 27MHz generated by this PLL
    pll0 : component pll 
        port map (
            refclk => i_clk_50,
            rst => not(i_rst_n),
            outclk_0 => s_clk_27,
            locked => s_rst_n
        );

    -- Configures the ADV7513 for 480p
    I2C_HDMI_Config0 : component I2C_HDMI_Config 
        port map (
            iCLK => i_clk_50,
            iRST_N => i_rst_n,
            I2C_SCLK => io_hdmi_i2c_scl,
            I2C_SDAT => io_hdmi_i2c_sda,
            HDMI_TX_INT => i_hdmi_tx_int
        );
    
    
    hdmi_controler : entity work.hdmi_controler
    generic map (
        H_RES => 720,
        V_RES => 480
    )
    port map (
        i_clk   => s_clk_27,
        i_rst_n => s_rst_n,
		  -- Sorties coordonnées
        o_x => s_scan_x,
        o_y => s_scan_y,  
        o_hdmi_tx_clk  => o_hdmi_tx_clk,
        o_hdmi_tx_de => s_de,
        o_hdmi_tx_hs   => o_hdmi_tx_hs,
        o_hdmi_tx_vs   => o_hdmi_tx_vs
    );
	 
	 -- Connexion de la sortie DE
    o_hdmi_tx_de <= s_de;
	
-- ========================================================================
    -- INSTANCIATION DES ENCODEURS 
    -- ========================================================================
    
    -- Encodeur Gauche (Axe X)
    inst_encoder_x : entity work.gestion_encodeur
    generic map (
        C_MAX_VAL   => h_res,    -- 720
        C_START_POS => h_res / 2 -- 360
    )
    port map (
        i_clk   => i_clk_50,
        i_rst_n => s_rst_n,
        i_a     => i_left_ch_a,
        i_b     => i_left_ch_b,
        o_val   => s_pos_x
    );

    -- Encodeur Droit (Axe Y)
    inst_encoder_y : entity work.gestion_encodeur
    generic map (
        C_MAX_VAL   => v_res,    -- 480
        C_START_POS => v_res / 2 -- 240
    )
    port map (
        i_clk   => i_clk_50,
        i_rst_n => s_rst_n,
        i_a     => i_right_ch_a,
        i_b     => i_right_ch_b,
        o_val   => s_pos_y
    );

	 -- ========================================================================
    -- AFFICHAGE (Carre Blanc sur Fond Bleu)
    -- ========================================================================
    -- AFFICHAGE
    process(s_clk_27) -- Utilise l'horloge HDMI, c'est plus propre que la liste de sensibilité
    begin
        if rising_edge(s_clk_27) then
            if s_de = '1' then
                -- Priorité au curseur (optionnel, pour voir où on est)
                if (to_integer(s_scan_x) >= s_pos_x and to_integer(s_scan_x) < s_pos_x + 4) and
                   (to_integer(s_scan_y) >= s_pos_y and to_integer(s_scan_y) < s_pos_y + 4) then
                    o_hdmi_tx_d <= x"00FF00"; -- Curseur Rouge
                
                -- Sinon, on affiche ce qu'il y a en mémoire
                elsif s_pixel_data(0) = '1' then
                    o_hdmi_tx_d <= x"000000"; 
                else
                    o_hdmi_tx_d <= x"00FF00"; 
                end if;
            else
                o_hdmi_tx_d <= (others => '0');
            end if;
        end if;
    end process;
	 
    -- Processus d'écriture dans la DPRAM via le port A
    process(i_left_pb, s_pos_x, s_pos_y)
    begin
         s_we_a   <= '1';
         s_data_a <= "1"; -- Vecteur de 1 bit à '1'
         s_addr_a <= s_pos_y * h_res + s_pos_x;

    end process;
	 
	-- DPRAM Instantiation
    inst_framebuffer : entity work.dpram
    generic map (
        mem_size   => h_res * v_res,
        data_width => 1  -- CORRECTION IMPORTANTE : 1 bit de large
    ) -- PAS DE POINT VIRGULE ICI !
    port map (    
        i_clk_a  => i_clk_50, -- Utilise i_clk_50 pour l'écriture (synchro avec encodeurs)
        i_clk_b  => s_clk_27, -- Utilise s_clk_27 pour la lecture (synchro avec HDMI)

        i_data_a => s_data_a,
        i_data_b => "0",      -- Vecteur de 1 bit
        i_addr_a => s_addr_a,
        i_addr_b => to_integer(s_scan_y) * h_res + to_integer(s_scan_x),
        i_we_a   => s_we_a,
        i_we_b   => '0',
        o_q_a    => open,
        o_q_b    => s_pixel_data
    );
	 
end architecture rtl;